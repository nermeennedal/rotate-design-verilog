module XOR(output reg [31:0] F,input [31:0] A ,input [31:0] B);
	always @(*) begin
	 F[0] = (A[0] & ~B[0]) | (~A[0] & B[0]);
	 F[1] = (A[1] & ~B[1]) | (~A[1] & B[1]);
	 F[2] = (A[2] & ~B[2]) | (~A[2] & B[2]);
	 F[3] = (A[3] & ~B[3]) | (~A[3] & B[3]);
	 F[4] = (A[4] & ~B[4]) | (~A[4] & B[4]);
	 F[5] = (A[5] & ~B[5]) | (~A[5] & B[5]);
	 F[6] = (A[6] & ~B[6]) | (~A[6] & B[6]);
	 F[7] = (A[7] & ~B[7]) | (~A[7] & B[7]);
	 F[8] = (A[8] & ~B[8]) | (~A[8] & B[8]);
	 F[9] = (A[9] & ~B[9]) | (~A[9] & B[9]);
	 F[10] = (A[10] & ~B[10]) | (~A[10] & B[10]);
	 F[11] = (A[11] & ~B[11]) | (~A[11] & B[11]);
	 F[12] = (A[12] & ~B[12]) | (~A[12] & B[12]);
	 F[13] = (A[13] & ~B[13]) | (~A[13] & B[13]);
	 F[14] = (A[14] & ~B[14]) | (~A[14] & B[14]);
	 F[15] = (A[15] & ~B[15]) | (~A[15] & B[15]);
	 F[16] = (A[16] & ~B[16]) | (~A[16] & B[16]);
	 F[17] = (A[17] & ~B[17]) | (~A[17] & B[17]);
	 F[18] = (A[18] & ~B[18]) | (~A[18] & B[18]);
	 F[19] = (A[19] & ~B[19]) | (~A[19] & B[19]);
	 F[20] = (A[20] & ~B[20]) | (~A[20] & B[20]);
	 F[21] = (A[21] & ~B[21]) | (~A[21] & B[21]);
	 F[22] = (A[22] & ~B[22]) | (~A[22] & B[22]);
	 F[23] = (A[23] & ~B[23]) | (~A[23] & B[23]);
	 F[24] = (A[24] & ~B[24]) | (~A[24] & B[24]);
	 F[25] = (A[25] & ~B[25]) | (~A[25] & B[25]);
	 F[26] = (A[26] & ~B[26]) | (~A[26] & B[26]);
	 F[27] = (A[27] & ~B[27]) | (~A[27] & B[27]);
	 F[28] = (A[28] & ~B[28]) | (~A[28] & B[28]);
	 F[29] = (A[29] & ~B[29]) | (~A[29] & B[29]);
	 F[30] = (A[30] & ~B[30]) | (~A[30] & B[30]);
	 F[31] = (A[31] & ~B[31]) | (~A[31] & B[31]);
 	end

endmodule
 
